`timescale 1ns/1ns
module Instruction_Memory (Addr, Data);
  
  input [31:0] Addr;
  
  output reg [31:0] Data;
  
  always @(Addr) begin
    case(Addr)
      0:   Data = 32'b1110_00_1_1101_0_0000_0000_000000010100; //1
      4:   Data = 32'b1110_00_1_1101_0_0000_0001_101000000001; //2
      8:   Data = 32'b1110_00_1_1101_0_0000_0010_000100000011; //3
      12:  Data = 32'b1110_00_0_0100_1_0010_0011_000000000010; //4
      16:  Data = 32'b1110_00_0_0101_0_0000_0100_000000000000; //5
      20:  Data = 32'b1110_00_0_0010_0_0100_0101_000100000100; //6
      24:  Data = 32'b1110_00_0_0110_0_0000_0110_000010100000; //7
      28:  Data = 32'b1110_00_0_1100_0_0101_0111_000101000010; //8
      32:  Data = 32'b1110_00_0_0000_0_0111_1000_000000000011;
      36:  Data = 32'b1110_00_0_1111_0_0000_1001_000000000110;
      40:  Data = 32'b1110_00_0_0001_0_0100_1010_000000000101;
      44:  Data = 32'b1110_00_0_1010_1_1000_0000_000000000110;
      48:  Data = 32'b0001_00_0_0100_0_0001_0001_000000000001;
      52:  Data = 32'b1110_00_0_1000_1_1001_0000_000000001000;
      56:  Data = 32'b0000_00_0_0100_0_0010_0010_000000000010;
      60:  Data = 32'b1110_00_1_1101_0_0000_0000_101100000001;
      64:  Data = 32'b1110_01_0_0100_0_0000_0001_000000000000;
      68:  Data = 32'b1110_01_0_0100_1_0000_1011_000000000000;
      72:  Data = 32'b1110_01_0_0100_0_0000_0010_000000000100;
      76:  Data = 32'b1110_01_0_0100_0_0000_0011_000000001000;
      80:  Data = 32'b1110_01_0_0100_0_0000_0100_000000001101;
      84:  Data = 32'b1110_01_0_0100_0_0000_0101_000000010000;
      88:  Data = 32'b1110_01_0_0100_0_0000_0110_000000010100;
      92:  Data = 32'b1110_01_0_0100_1_0000_1010_000000000100;
      96:  Data = 32'b1110_01_0_0100_0_0000_0111_000000011000;
      100: Data = 32'b1110_00_1_1101_0_0000_0001_000000000100;
      104: Data = 32'b1110_00_1_1101_0_0000_0010_000000000000;
      108: Data = 32'b1110_00_1_1101_0_0000_0011_000000000000;
      112: Data = 32'b1110_00_0_0100_0_0000_0100_000100000011;
      116: Data = 32'b1110_01_0_0100_1_0100_0101_000000000000;
      120: Data = 32'b1110_01_0_0100_1_0100_0110_000000000100;
      124: Data = 32'b1110_00_0_1010_1_0101_0000_000000000110;
      128: Data = 32'b1100_01_0_0100_0_0100_0110_000000000000;
      132: Data = 32'b1100_01_0_0100_0_0100_0101_000000000100;
      136: Data = 32'b1110_00_1_0100_0_0011_0011_000000000001;
      140: Data = 32'b1110_00_1_1010_1_0011_0000_000000000011;
      144: Data = 32'b1011_10_1_0_111111111111111111110111;
      148: Data = 32'b1110_00_1_0100_0_0010_0010_000000000001;
      152: Data = 32'b1110_00_0_1010_1_0010_0000_000000000001;
      156: Data = 32'b1011_10_1_0_111111111111111111110011;
      160: Data = 32'b1110_01_0_0100_1_0000_0001_000000000000;
      164: Data = 32'b1110_01_0_0100_1_0000_0010_000000000100;
      168: Data = 32'b1110_01_0_0100_1_0000_0011_000000001000;
      172: Data = 32'b1110_01_0_0100_1_0000_0100_000000001100;
      176: Data = 32'b1110_01_0_0100_1_0000_0101_000000010000;
      180: Data = 32'b1110_01_0_0100_1_0000_0110_000000010100;
      184: Data = 32'b1110_10_1_0_111111111111111111111111;
      default: Data = 32'd0;
    endcase
  end
  
endmodule



module IM_TB();
  
  reg [31:0] Addr;
  
  wire [31:0] Data;
  
  Instruction_Memory uut(Addr, Data);
  
  
  initial begin
    Addr = 2;
    #20;
    Addr = 4;
    #20;
    Addr = 6;
    #20;
    Addr = 7;
    #20; 
  end
  
endmodule
  
